module and2x1 (out,in1,in2);
input in1,in2;
output out;

assign out = in1 & in2 ;

endmodule
