module not1x1 (out,in)
input in;
output out;

assign out = ~in;

endmodule
